
LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY gerador_de_paridade IS
port(	a: in std_logic;
	b: in std_logic;
	c: in std_logic;
	P: out std_logic
);

END gerador_de_paridade;

ARCHITECTURE logica OF gerador_de_paridade IS
	
BEGIN
	P <= a XOR b XOR c;
	
END logica;
